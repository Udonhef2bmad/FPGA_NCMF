LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;

ENTITY toplevel IS 
END ENTITY;

ARCHITECTURE RTL OF toplevel IS

BEGIN

END ARCHITECTURE;