COUNTER_inst : COUNTER PORT MAP (
		clock	 => clock_sig,
		updown	 => updown_sig,
		q	 => q_sig
	);
